[DMP3098L]
*DIODES_INC_SPICE_MODEL DMP3098L 
*SIMULATOR=SIMETRIX
*ORIGIN=DZSL_DPG_SU
*DATE=11Dec2012
*VERSION=1

.SUBCKT DMP3098L   10 20 30
M1 1 2 3 3  Pmod1
RD 10 1 Rmod1 27E-3
RS 23 3 Rmod1 27E-3
RG 20 22 5
RIN 20 23 2E11
RDS 10 23 2E9
CGS 2 3 100E-12 
EGD 12 0 1 2 1
REGD 12 0 1
VFB 14 0 0 
FFB 1 2 VFB 1 
CGD 13 14 400E-12 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 10 23 DSUB
EL 2 22 1 3 .003
RL 30 23 3
LS  30 23 2E-9
.MODEL Pmod1 PMOS (LEVEL=3 VTO=-2.1 TOX=6E-8 NSUB=5E+16 KP=9 NFS=1E11 IS=1E-15 N=10)
.MODEL DCGD D (CJO = 350E-12  VJ = 0.45  M = 0.33)
.MODEL DSUB D (IS=2.5E-13 N=1 RS=0.018 BV=33 CJO=94E-12 VJ=0.45 M=0.33 TT=3E-9)
.MODEL DLIM D (IS=100U N=1)
.MODEL Rmod1 RES (TC1=.5e-3 TC2=3E-6)
.ENDS