**********************************
**********************************
**
** Littelfuse, Inc
** TVS Diode SPICE Models
** SMBJxxxCA
**
** Jifeng Z.
** Wuxi Technical Center
**
** A 01/06/2012
** MODEL FORMAT: SPICE3
**
**********************************
**********************************
.SUBCKT SMBJ24CA   1  2
*       TERMINALS: T1 T2
Done    1          3  Dtvs
Dtwo    2          3  Dtvs
Rleak   1          2  48meg
.MODEL  Dtvs       D  (IS=1.0e-5 RS=0.0983 N=1.5 IBV=1m BV=26.97 CJO=900p)
.ENDS
