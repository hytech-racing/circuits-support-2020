*---------- DMP3099L Spice Model ----------
.SUBCKT DMP3099L D G S
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006
RD 10 1 0.02942
RS 30 3 0.001
RG 20 2 10.27
CGS 2 3 5.366E-010
EGD 12 30 2 1 1
VFB 14 30 0
FFB 2 1 VFB 1
CGD 13 14 4.4E-010
R1 13 30 1
D1 13 12 DLIM
DDG 14 15 DCGD
R2 12 15 1
D2 30 15 DLIM
DSD 10 3 DSUB
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 TOX = 6E-008 NSUB = 1E+016 KP = 8.769 KAPPA = 19.32 VTO = -1.917
.MODEL DCGD D CJO = 2.502E-010 VJ = 0.8 M = 0.6
.MODEL DSUB D IS = 4.949E-009 N = 1.628 RS = 0.02235 BV = 33 CJO = 5.295E-011 VJ = 0.8 M = 0.6
.MODEL DLIM D IS = 0.0001
.ENDS
*Diodes DMP3099L Spice Model v1.0M Last Revised 2017/12/7